library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity IM is
    port (
		    rst  : in std_logic;
        addr : in  std_logic_vector(31 downto 0);
        data : out std_logic_vector(31 downto 0)
    );
end IM;

architecture behavioral of IM is
    type memoria_rom is array (0 to 63) of std_logic_vector (31 downto 0);
    signal ROM : memoria_rom := (
"10000010000100000010000000000101", --mov  5, %g1
"10100000000100000011111111111000", --mov  -8, %l0
"10100010000100000010000000000100", --mov  4, %l1
"10110001001010000110000000000010", --sll %g1, 2, %i0
"10110011001101000110000000000001", --srl %l1, 1, %i1
"10000001111010000010000000000000",--restore %g0,0,%g0
"10100000000000000110000000000011", --add %g1,3,%l0
"10000001111000000010000000000000",--save %g0,0,%g0
"10000000101000000010000000000100", -- subcc %g0,4,%g0
"00000000000000000000000000000000",
"10000100010000000000000000000001", -- addx %g0,%g1, %g2
"10010000000100000000000000010000", -- mov %l0, %o0
"00000001000000000000000000000000", --nop
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
--"00000000000000000000000000000000",
--"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000" -- Fila con datos 56 a 63
    );
begin
	process(rst, addr)
	begin
	 if (rst = '1') then
			data <= "00000000000000000000000000000000";
		else
			data <= ROM(conv_integer(addr));
	 end if;
	end process;
end behavioral;




--from random import randint

--n = 64

--for i in xrange(n):
   -- x = randint(0, 1<<32)
    --num = str(bin(x))[2:]
    --num = (32 - len(num)) * '0' + num
    --print "\"" + num + "\","
